parameter   FT600_CLK_PERIOD = 4,
parameter   MAIN_CLK_PERIOD = 3