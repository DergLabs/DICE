parameter   DDR_CLK_PERIOD = 5000,
parameter   MAIN_CLK_PERIOD = 10000